

`include "uvm_macros.svh"
package uart_responder_tests_pkg;
	import uvm_pkg::*;
	import uart_responder_env_pkg::*;
	
	`include "uart_responder_test_base.svh"
	
endpackage
