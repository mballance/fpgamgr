
`include "uvm_macros.svh"

package uart_responder_env_pkg;
	import uvm_pkg::*;

	`include "uart_responder_env.svh"
	
endpackage
